// basic module to interface with adxl345 accelerometer. This will initialize
// the device and place it in FIFO mode. The resulting the stream will be
// collected by the SPI master peripheral. The resulting stream will contain the
// x, y, z data of the accelerometer
`timescale 1ns / 1ps
`default_nettype none

module adxl345 ();
    // TODO
endmodule

`default_nettype wire
