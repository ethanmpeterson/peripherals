`timescale 1ns / 1ps
`default_nettype none

module mdio_master;
endmodule

`default_nettype wire
