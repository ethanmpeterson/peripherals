`default_nettype none
`timescale 1ns / 1ps

interface axis_interface ();

endinterface // mdio_interface

`default_nettype wire
