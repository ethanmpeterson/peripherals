`timescale 1ns / 1ps
`default_nettype none

module dp83848x;
endmodule

`default_nettype wire