`timescale 1ns / 1ps
`default_nettype none

module adxl345_bfm (
    spi_interface.slave spi_bus,
);

endmodule

`default_nettype wire
