`default_nettype none
`timescale 1ns / 1ps

module udp_checksum_gen_wrapper (
);

endmodule

`default_nettype wire
